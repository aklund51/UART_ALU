`timescale 1ns / 1ps

package config_pkg;

// define structs and enums needed for design

endpackage
