module uart_alu (
    input clk_12mhz_i,
    input reset_unsafe_i
);
    
endmodule
