package config_pkg;

// define structs and enums needed for design

endpackage
